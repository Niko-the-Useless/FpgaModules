module greaterThan
(
	input [3:0] i_a,
	input [3:0] i_b,
	output o_ab
);
	assign o_ab=(i_a>i_b);
endmodule
